CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 1532 489
9961490 0
0
6 Title:
5 Name:
0
0
0
9
7 Ground~
168 421 332 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
4212 0 0
2
5.89879e-315 0
0
11 Multimeter~
205 527 24 0 21 21
0 3 7 8 4 0 0 0 0 0
32 52 51 48 46 52 109 86 0 0
0 82
0
0 0 16464 0
8 100.0Meg
-28 -19 28 -11
3 MM2
-11 -29 10 -21
0
0
11 %D %1 %4 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
1 R
4720 0 0
2
5.89879e-315 0
0
11 Multimeter~
205 343 31 0 21 21
0 5 9 10 3 0 0 0 0 0
32 49 57 46 50 55 32 86 0 0
0 82
0
0 0 16464 0
8 100.0Meg
-28 -19 28 -11
3 MM1
-11 -29 10 -21
0
0
11 %D %1 %4 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
1 R
5551 0 0
2
5.89879e-315 0
0
11 Multimeter~
205 531 158 0 21 21
0 3 11 12 6 0 0 0 0 0
32 49 56 46 51 53 109 65 0 0
0 86
0
0 0 16464 270
6 1.000u
-21 -19 21 -11
3 MM0
-11 -29 10 -21
0
0
28 R1%D %1 %2 %V
%D %2 %4 DC 0
0
0
0
9

0 1 2 3 4 1 2 3 4 0
86 0 0 0 1 0 0 0
1 V
6986 0 0
2
5.89879e-315 0
0
6 Diode~
219 407 171 0 2 5
0 6 2
0
0 0 848 270
5 DIODE
11 0 46 8
2 D1
22 -10 36 -2
0
0
11 %D %1 %2 %M
0
0
9 DOIODE0.4
5

0 -54 -44 -54 -44 0
68 0 0 0 1 0 0 0
1 D
8745 0 0
2
5.89879e-315 0
0
8 Battery~
219 656 217 0 2 5
0 4 2
0
0 0 880 0
3 0.3
12 -2 33 6
2 Ge
16 -12 30 -4
0
0
14 %D %1 %2 DC %V
0
0
0
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
1 V
9592 0 0
2
5.89879e-315 0
0
8 Battery~
219 244 195 0 2 5
0 5 2
0
0 0 880 0
3 20V
12 -2 33 6
2 V1
15 -12 29 -4
0
0
14 %D %1 %2 DC %V
0
0
0
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
1 V
8748 0 0
2
5.89879e-315 0
0
9 Resistor~
219 537 102 0 2 5
0 3 4
0
0 0 880 0
9 0.47k Ohm
-31 -14 32 -6
2 R2
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
7168 0 0
2
5.89879e-315 0
0
9 Resistor~
219 342 102 0 2 5
0 5 3
0
0 0 880 0
6 1k Ohm
-21 -14 21 -6
2 R1
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
631 0 0
2
5.89879e-315 0
0
12
4 0 3 0 0 4096 0 3 0 0 11 2
368 54
368 102
2 0 2 0 0 4096 0 5 0 0 5 2
407 181
407 277
0 1 2 0 0 0 0 0 1 5 0 4
406 277
406 318
421 318
421 326
4 0 4 0 0 4096 0 2 0 0 6 4
552 47
552 94
568 94
568 102
2 2 2 0 0 8320 0 6 7 0 0 4
656 228
656 277
244 277
244 206
2 1 4 0 0 8320 0 8 6 0 0 3
555 102
656 102
656 204
1 0 3 0 0 4096 0 2 0 0 11 4
502 47
502 97
503 97
503 102
1 0 5 0 0 4096 0 3 0 0 12 2
318 54
318 102
1 0 3 0 0 4096 0 4 0 0 11 3
515 140
422 140
422 102
4 1 6 0 0 8320 0 4 5 0 0 6
515 190
515 146
394 146
394 153
407 153
407 161
2 1 3 0 0 4224 0 9 8 0 0 2
360 102
519 102
1 1 5 0 0 4224 0 7 9 0 0 3
244 182
244 102
324 102
0
0
2049 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
