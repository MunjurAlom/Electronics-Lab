CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 1532 489
9961490 0
0
6 Title:
5 Name:
0
0
0
9
7 Ground~
168 398 420 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
9196 0 0
2
43496.8 0
0
8 Battery~
219 271 197 0 2 5
0 3 2
0
0 0 880 0
3 10V
12 -2 33 6
2 V1
16 -12 30 -4
0
0
14 %D %1 %2 DC %V
0
0
0
5

0 1 2 1 2 0
86 0 0 0 0 0 0 0
1 V
3857 0 0
2
43496.8 0
0
11 Multimeter~
205 791 223 0 21 21
0 4 8 9 2 0 0 0 0 0
32 54 46 50 50 50 32 86 0 0
0 82
0
0 0 16464 0
8 100.0Meg
-28 -19 28 -11
3 MM1
-11 -29 10 -21
0
0
11 %D %1 %4 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 0 0 0 0
1 R
7125 0 0
2
43496.8 0
0
11 Multimeter~
205 309 82 0 21 21
0 3 10 11 5 0 0 0 0 0
32 49 46 53 53 53 109 65 0 0
0 86
0
0 0 16464 0
6 1.000u
-21 -19 21 -11
3 MM0
-11 -29 10 -21
0
0
28 R1%D %1 %2 %V
%D %2 %4 DC 0
0
0
0
9

0 1 2 3 4 1 2 3 4 0
86 0 0 0 0 0 0 0
1 V
3641 0 0
2
43496.8 0
0
6 Diode~
219 374 252 0 2 5
0 3 7
0
0 0 848 0
5 DIODE
-18 -18 17 -10
2 D2
-7 -28 7 -20
0
0
11 %D %1 %2 %M
0
0
9 DOIODE0.4
5

0 -54 -44 -54 -44 0
68 0 0 0 0 0 0 0
1 D
9821 0 0
2
43496.8 0
0
6 Diode~
219 387 127 0 2 5
0 5 6
0
0 0 848 0
5 DIODE
-18 -18 17 -10
2 D1
-7 -28 7 -20
0
0
11 %D %1 %2 %M
0
0
9 DOIODE0.4
5

0 -54 -44 -54 -44 0
68 0 0 0 0 0 0 0
1 D
3187 0 0
2
43496.8 0
0
9 Resistor~
219 669 283 0 3 5
0 2 4 -1
0
0 0 880 90
6 2k Ohm
-6 0 36 8
2 R3
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 0 0 0 0
1 R
762 0 0
2
43496.8 0
0
9 Resistor~
219 515 240 0 2 5
0 7 4
0
0 0 880 0
6 2k Ohm
-20 -14 22 -6
2 R2
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 0 0 0 0
1 R
39 0 0
2
43496.8 0
0
9 Resistor~
219 517 170 0 2 5
0 6 4
0
0 0 880 0
6 2k Ohm
-21 -14 21 -6
2 R1
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 0 0 0 0
1 R
9450 0 0
2
43496.8 0
0
11
1 0 3 0 0 4096 0 4 0 0 7 2
284 105
284 168
1 0 2 0 0 4096 0 1 0 0 5 2
398 414
398 368
4 0 2 0 0 8192 0 3 0 0 5 3
816 246
816 323
669 323
1 0 4 0 0 8192 0 3 0 0 8 3
766 246
766 250
669 250
2 1 2 0 0 8320 0 2 7 0 0 4
271 208
271 368
669 368
669 301
4 1 5 0 0 8320 0 4 6 0 0 3
334 105
334 127
377 127
1 1 3 0 0 8336 0 2 5 0 0 5
271 184
271 168
356 168
356 252
364 252
0 2 4 0 0 4224 0 0 7 10 0 3
543 203
669 203
669 265
1 2 6 0 0 4224 0 9 6 0 0 4
499 170
405 170
405 127
397 127
2 2 4 0 0 0 0 8 9 0 0 4
533 240
543 240
543 170
535 170
2 1 7 0 0 4224 0 5 8 0 0 4
384 252
489 252
489 240
497 240
0
0
2049 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
