CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
176 80 1364 717
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.499215 0.500000
344 176 1532 493
9961490 0
0
6 Title:
5 Name:
0
0
0
8
11 Multimeter~
205 372 183 0 21 21
0 3 7 8 4 0 0 0 0 0
32 54 46 57 53 50 109 65 0 0
0 86
0
0 0 16464 180
6 1.000u
-21 -19 21 -11
3 MM5
-11 -29 10 -21
0
0
28 R1%D %1 %2 %V
%D %2 %4 DC 0
0
0
0
9

0 1 2 3 4 1 2 3 4 0
86 0 0 0 0 0 0 0
1 V
5130 0 0
2
43475.8 0
0
7 Ground~
168 782 368 0 1 3
0 2
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
391 0 0
2
43475.8 0
0
8 Battery~
219 738 222 0 2 5
0 2 5
0
0 0 880 270
2 4V
-8 -20 6 -12
2 E2
-7 -30 7 -22
0
0
14 %D %1 %2 DC %V
0
0
0
5

0 1 2 1 2 0
86 0 0 0 0 0 0 0
1 V
3124 0 0
2
43475.8 0
0
7 Ground~
168 297 364 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
3421 0 0
2
43475.8 0
0
6 Diode~
219 557 263 0 2 5
0 5 6
0
0 0 848 180
5 DIODE
-18 -18 17 -10
2 D2
-7 -28 7 -20
0
0
11 %D %1 %2 %M
0
0
9 DOIODE0.4
5

0 -54 -44 -54 -44 0
68 0 0 0 0 0 0 0
1 D
8157 0 0
2
43475.8 0
0
6 Diode~
219 549 164 0 2 5
0 6 5
0
0 0 848 0
5 DIODE
-18 -18 17 -10
2 D1
-7 -28 7 -20
0
0
11 %D %1 %2 %M
0
0
9 DOIODE0.4
5

0 -54 -44 -54 -44 0
68 0 0 0 0 0 0 0
1 D
5572 0 0
2
43475.8 0
0
8 Battery~
219 301 215 0 2 5
0 2 4
0
0 0 880 90
3 20V
-10 -21 11 -13
2 E1
-7 -31 7 -23
0
0
14 %D %1 %2 DC %V
0
0
0
5

0 1 2 1 2 0
86 0 0 0 0 0 0 0
1 V
8901 0 0
2
43475.8 0
0
9 Resistor~
219 435 212 0 2 5
0 3 6
0
0 0 880 0
8 2.2k Ohm
-19 -17 37 -9
2 R1
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 0 0 0 0
1 R
7361 0 0
2
43475.8 0
0
8
1 1 3 0 0 8320 0 8 1 0 0 5
417 212
413 212
413 170
395 170
395 174
4 2 4 0 0 12432 0 1 7 0 0 5
345 174
345 172
327 172
327 212
315 212
1 1 2 0 0 8320 0 3 2 0 0 3
749 220
782 220
782 362
1 1 2 0 0 0 0 7 4 0 0 5
291 212
279 212
279 350
297 350
297 358
2 0 5 0 0 4096 0 3 0 0 6 2
725 220
635 220
2 1 5 0 0 8320 0 6 5 0 0 4
559 164
635 164
635 263
567 263
2 0 6 0 0 4096 0 8 0 0 8 2
453 212
493 212
2 1 6 0 0 8320 0 5 6 0 0 4
547 263
493 263
493 164
539 164
0
0
2049 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
