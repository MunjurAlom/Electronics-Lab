CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
176 80 1364 717
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 1532 494
9961490 0
0
6 Title:
5 Name:
0
0
0
9
11 Multimeter~
205 817 188 0 21 21
0 4 7 8 2 0 0 0 0 0
32 54 52 56 46 52 117 86 0 0
0 82
0
0 0 16464 270
8 100.0Meg
-28 -19 28 -11
3 MM2
-11 -29 10 -21
0
0
11 %D %1 %4 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 0 0 0 0
1 R
7361 0 0
2
43468.9 0
0
11 Multimeter~
205 659 42 0 21 21
0 5 9 10 4 0 0 0 0 0
32 49 49 46 53 56 32 86 0 0
0 82
0
0 0 16464 0
8 100.0Meg
-28 -19 28 -11
3 MM1
-11 -29 10 -21
0
0
11 %D %1 %4 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 0 0 0 0
1 R
4747 0 0
2
43468.9 0
0
11 Multimeter~
205 474 56 0 21 21
0 3 11 12 5 0 0 0 0 0
32 49 49 53 46 56 110 65 0 0
0 86
0
0 0 16464 0
6 1.000u
-21 -19 21 -11
3 MM0
-11 -29 10 -21
0
0
28 R1%D %1 %2 %V
%D %2 %4 DC 0
0
0
0
9

0 1 2 3 4 1 2 3 4 0
86 0 0 0 0 0 0 0
1 V
972 0 0
2
43468.9 0
0
6 Diode~
219 640 127 0 2 5
0 4 5
0
0 0 848 180
5 DIODE
-18 -18 17 -10
2 D2
-7 -28 7 -20
0
0
11 %D %1 %2 %M
0
0
9 DOIODE0.4
5

0 -54 -44 -54 -44 0
68 0 0 0 0 0 0 0
1 D
3472 0 0
2
43468.9 0
0
6 Diode~
219 488 126 0 2 5
0 6 3
0
0 0 848 0
5 DIODE
-18 -18 17 -10
2 D1
-7 -28 7 -20
0
0
11 %D %1 %2 %M
0
0
9 DOIODE0.4
5

0 -54 -44 -54 -44 0
68 0 0 0 0 0 0 0
1 D
9998 0 0
2
43468.9 0
0
7 Ground~
168 646 314 0 1 3
0 2
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
3536 0 0
2
43468.9 0
0
7 Ground~
168 411 320 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
4597 0 0
2
43468.9 0
0
8 Battery~
219 392 165 0 2 5
0 6 2
0
0 0 880 0
3 12V
12 -2 33 6
2 V1
16 -12 30 -4
0
0
14 %D %1 %2 DC %V
0
0
0
5

0 1 2 1 2 0
86 0 0 0 0 0 0 0
1 V
3835 0 0
2
43468.9 0
0
9 Resistor~
219 718 188 0 3 5
0 2 4 -1
0
0 0 880 90
8 5.6k Ohm
11 -1 67 7
2 R1
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 0 0 0 0
1 R
3670 0 0
2
43468.9 0
0
10
2 1 3 0 0 12416 0 5 3 0 0 5
498 126
516 126
516 92
449 92
449 79
4 0 2 0 0 8320 0 1 0 0 6 3
801 220
801 270
718 270
0 1 4 0 0 4224 0 0 1 4 0 4
717 127
794 127
794 170
801 170
4 0 4 0 0 0 0 2 0 0 9 3
684 65
717 65
717 127
1 0 5 0 0 8192 0 2 0 0 7 3
634 65
606 65
606 127
1 1 2 0 0 0 0 6 9 0 0 4
646 308
646 270
718 270
718 206
4 2 5 0 0 4240 0 3 4 0 0 4
499 79
592 79
592 127
630 127
2 1 2 0 0 0 0 8 7 0 0 6
392 176
392 225
361 225
361 252
411 252
411 314
1 2 4 0 0 0 0 4 9 0 0 3
650 127
718 127
718 170
1 1 6 0 0 8320 0 8 5 0 0 3
392 152
392 126
478 126
0
0
2049 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
