CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 1532 489
9961490 0
0
6 Title:
5 Name:
0
0
0
10
11 Multimeter~
205 755 297 0 21 21
0 3 8 9 4 0 0 0 0 0
32 52 46 53 54 56 32 86 0 0
0 82
0
0 0 16464 270
8 100.0Meg
-28 -19 28 -11
3 MM3
-11 -29 10 -21
0
0
11 %D %1 %4 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 0 0 0 0
1 R
3409 0 0
2
43539 0
0
11 Multimeter~
205 924 352 0 21 21
0 3 10 11 2 0 0 0 0 0
45 52 51 50 46 50 109 86 0 0
0 82
0
0 0 16464 270
8 100.0Meg
-28 -19 28 -11
3 MM2
-11 -29 10 -21
0
0
11 %D %1 %4 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 0 0 0 0
1 R
3951 0 0
2
43539 0
0
11 Multimeter~
205 631 180 0 21 21
0 5 12 13 3 0 0 0 0 0
32 50 46 48 55 54 109 65 0 0
0 86
0
0 0 16464 0
6 1.000u
-21 -19 21 -11
3 MM1
-11 -29 10 -21
0
0
28 R1%D %1 %2 %V
%D %2 %4 DC 0
0
0
0
9

0 1 2 3 4 1 2 3 4 0
86 0 0 0 0 0 0 0
1 V
8885 0 0
2
43539 0
0
11 Multimeter~
205 420 147 0 21 21
0 7 14 15 6 0 0 0 0 0
32 57 46 55 53 56 32 86 0 0
0 82
0
0 0 16464 0
8 100.0Meg
-28 -19 28 -11
3 MM0
-11 -29 10 -21
0
0
11 %D %1 %4 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 0 0 0 0
1 R
3780 0 0
2
43539 0
0
7 Ground~
168 332 510 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
9265 0 0
2
43539 0
0
8 Battery~
219 691 417 0 2 5
0 2 4
0
0 0 880 180
2 5V
14 -2 28 6
2 V2
15 -12 29 -4
0
0
14 %D %1 %2 DC %V
0
0
0
5

0 1 2 1 2 0
86 0 0 0 0 0 0 0
1 V
9442 0 0
2
43539 0
0
6 Diode~
219 547 229 0 2 5
0 6 5
0
0 0 848 0
5 DIODE
-18 -18 17 -10
2 D1
-7 -28 7 -20
0
0
11 %D %1 %2 %M
0
0
9 DOIODE0.4
5

0 -54 -44 -54 -44 0
68 0 0 0 0 0 0 0
1 D
9424 0 0
2
43539 0
0
8 Battery~
219 306 231 0 2 5
0 7 2
0
0 0 880 270
3 10V
-11 -20 10 -12
2 V1
-7 -30 7 -22
0
0
14 %D %1 %2 DC %V
0
0
0
5

0 1 2 1 2 0
86 0 0 0 0 0 0 0
1 V
9968 0 0
2
43539 0
0
9 Resistor~
219 689 307 0 2 5
0 4 3
0
0 0 880 90
4 2.2k
1 0 29 8
2 R2
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 0 0 0 0
1 R
9281 0 0
2
43539 0
0
9 Resistor~
219 422 229 0 2 5
0 7 6
0
0 0 880 0
4 4.7k
-14 -14 14 -6
2 R1
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 0 0 0 0
1 R
8464 0 0
2
43539 0
0
13
1 0 3 0 0 4240 0 2 0 0 8 5
908 334
775 334
775 234
687 234
687 233
1 0 3 0 0 0 0 1 0 0 8 4
739 279
694 279
694 280
689 280
0 4 2 0 0 4096 0 0 2 7 0 4
689 444
900 444
900 384
908 384
4 0 4 0 0 4096 0 1 0 0 5 2
739 329
689 329
1 2 4 0 0 4224 0 9 6 0 0 2
689 325
689 402
1 0 2 0 0 0 0 5 0 0 7 2
332 504
332 461
1 2 2 0 0 8320 0 6 8 0 0 5
689 426
689 461
225 461
225 229
293 229
4 2 3 0 0 0 0 3 9 0 0 4
656 203
656 233
689 233
689 289
2 1 5 0 0 4224 0 7 3 0 0 3
557 229
606 229
606 203
4 0 6 0 0 4096 0 4 0 0 12 2
445 170
445 229
1 0 7 0 0 4096 0 4 0 0 13 2
395 170
395 229
2 1 6 0 0 4224 0 10 7 0 0 2
440 229
537 229
1 1 7 0 0 4224 0 8 10 0 0 2
317 229
404 229
0
0
2049 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
