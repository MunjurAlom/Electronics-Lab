CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
176 80 1364 717
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 1532 494
9961490 0
0
6 Title:
5 Name:
0
0
0
8
11 Multimeter~
205 762 264 0 21 21
0 3 7 8 2 0 0 0 0 0
32 55 49 50 46 55 109 86 0 0
0 82
0
0 0 16464 0
8 100.0Meg
-28 -19 28 -11
3 MM2
-11 -29 10 -21
0
0
11 %D %1 %4 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 0 0 0 0
1 R
9466 0 0
2
43478.8 0
0
8 Battery~
219 663 409 0 2 5
0 6 2
0
0 0 880 0
3 10V
12 -2 33 6
1 E
19 -12 26 -4
0
0
14 %D %1 %2 DC %V
0
0
0
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
1 V
3266 0 0
2
5.89877e-315 0
0
6 Diode~
219 533 269 0 2 5
0 3 4
0
0 0 848 180
5 DIODE
-18 -18 17 -10
2 D2
-7 -28 7 -20
0
0
11 %D %1 %2 %M
0
0
9 DOIODE0.4
5

0 -54 -44 -54 -44 0
68 0 0 0 1 0 0 0
1 D
7693 0 0
2
5.89877e-315 0
0
8 Battery~
219 430 283 0 2 5
0 4 2
0
0 0 880 270
2 0V
-7 -20 7 -12
2 E2
-7 -30 7 -22
0
0
14 %D %1 %2 DC %V
0
0
0
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
1 V
3723 0 0
2
5.89877e-315 0
0
6 Diode~
219 531 202 0 2 5
0 3 5
0
0 0 848 180
5 DIODE
-18 -18 17 -10
2 D1
-7 -28 7 -20
0
0
11 %D %1 %2 %M
0
0
9 DOIODE0.4
5

0 -54 -44 -54 -44 0
68 0 0 0 1 0 0 0
1 D
3440 0 0
2
5.89877e-315 0
0
7 Ground~
168 472 476 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
6263 0 0
2
5.89877e-315 0
0
8 Battery~
219 425 222 0 2 5
0 5 2
0
0 0 880 0
3 10V
12 -2 33 6
2 E1
16 -12 30 -4
0
0
14 %D %1 %2 DC %V
0
0
0
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
1 V
4900 0 0
2
5.89877e-315 0
0
9 Resistor~
219 659 322 0 2 5
0 6 3
0
0 0 880 90
2 1k
8 0 22 8
1 R
11 -10 18 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
8783 0 0
2
5.89877e-315 0
0
10
4 0 2 0 0 4096 0 1 0 0 6 3
787 287
787 440
663 440
1 0 3 0 0 8192 0 1 0 0 3 3
737 287
737 291
659 291
0 2 3 0 0 4224 0 0 8 4 0 3
551 234
659 234
659 304
1 1 3 0 0 0 0 5 3 0 0 4
541 202
551 202
551 269
543 269
1 0 2 0 0 0 0 6 0 0 6 2
472 470
472 455
2 0 2 0 0 8320 0 2 0 0 8 4
663 420
663 455
404 455
404 281
1 2 4 0 0 4224 0 4 3 0 0 4
441 281
515 281
515 269
523 269
2 2 2 0 0 0 0 7 4 0 0 4
425 233
404 233
404 281
417 281
1 2 5 0 0 8320 0 7 5 0 0 5
425 209
425 198
513 198
513 202
521 202
1 1 6 0 0 12416 0 2 8 0 0 4
663 396
663 371
659 371
659 340
0
0
2049 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
