CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
176 80 1364 717
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 1532 494
9961490 0
0
6 Title:
5 Name:
0
0
0
6
6 Diode~
219 400 274 0 2 5
0 4 3
0
0 0 848 270
5 DIODE
11 0 46 8
2 D1
22 -10 36 -2
0
0
11 %D %1 %2 %M
0
0
9 DOIODE0.4
5

0 -54 -44 -54 -44 0
68 0 0 0 0 0 0 0
1 D
4747 0 0
2
43475.8 0
0
8 Battery~
219 264 334 0 2 5
0 4 2
0
0 0 880 0
3 12V
12 -2 33 6
2 V1
16 -12 30 -4
0
0
14 %D %1 %2 DC %V
0
0
0
5

0 1 2 1 2 0
86 0 0 0 0 0 0 0
1 V
972 0 0
2
43475.8 0
0
11 Multimeter~
205 598 389 0 21 21
0 3 5 6 2 0 0 0 0 0
32 49 49 46 55 48 32 86 0 0
0 82
0
0 0 16464 270
8 100.0Meg
-28 -19 28 -11
3 MM0
-11 -29 10 -21
0
0
11 %D %1 %4 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 0 0 0 0
1 R
3472 0 0
2
43475.8 0
0
7 Ground~
168 328 525 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
9998 0 0
2
43475.8 0
0
8 Battery~
219 467 273 0 2 5
0 4 3
0
0 0 880 0
3 0.3
12 -2 33 6
2 V2
16 -12 30 -4
0
0
14 %D %1 %2 DC %V
0
0
0
5

0 1 2 1 2 0
86 0 0 0 0 0 0 0
1 V
3536 0 0
2
43475.8 0
0
9 Resistor~
219 460 391 0 3 5
0 2 3 -1
0
0 0 880 90
4 2.2k
1 0 29 8
2 R1
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 0 0 0 0
1 R
4597 0 0
2
43475.8 0
0
8
1 0 3 0 0 4224 0 3 0 0 8 4
582 371
468 371
468 325
435 325
1 0 4 0 0 8192 0 5 0 0 3 4
467 260
467 249
400 249
400 256
1 1 4 0 0 8320 0 2 1 0 0 4
264 321
264 256
400 256
400 264
2 2 3 0 0 16 0 5 1 0 0 4
467 284
467 310
400 310
400 284
4 0 2 0 0 4096 0 3 0 0 7 2
582 421
460 421
0 1 2 0 0 0 0 0 4 7 0 2
328 462
328 519
2 1 2 0 0 8320 0 2 6 0 0 4
264 345
264 462
460 462
460 409
0 2 3 0 0 0 0 0 6 4 0 4
435 310
435 333
460 333
460 373
0
0
2049 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
