CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
176 80 1364 717
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.499215 0.500000
344 176 1532 493
9961490 0
0
6 Title:
5 Name:
0
0
0
7
11 Multimeter~
205 671 163 0 21 21
0 3 7 8 2 0 0 0 0 0
32 49 49 46 48 48 32 86 0 0
0 82
0
0 0 16464 270
8 100.0Meg
-28 -19 28 -11
3 MM1
-11 -29 10 -21
0
0
11 %D %1 %4 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 0 0 0 0
1 R
5130 0 0
2
43468.9 0
0
11 Multimeter~
205 282 145 0 21 21
0 5 9 10 4 0 0 0 0 0
32 49 46 57 54 52 109 65 0 0
0 86
0
0 0 16464 90
6 1.000u
-21 -19 21 -11
3 MM0
-11 -29 10 -21
0
0
28 R1%D %1 %2 %V
%D %2 %4 DC 0
0
0
0
9

0 1 2 3 4 1 2 3 4 0
86 0 0 0 0 0 0 0
1 V
391 0 0
2
43468.9 0
0
7 Ground~
168 373 281 0 1 3
0 11
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 512 0 0 0 0
3 GND
3124 0 0
2
43468.9 0
0
8 Battery~
219 441 109 0 2 5
0 6 3
0
0 0 880 90
3 0.3
-11 -21 10 -13
2 V2
-8 -31 6 -23
0
0
14 %D %1 %2 DC %V
0
0
0
5

0 1 2 1 2 0
86 0 0 0 0 0 0 0
1 V
3421 0 0
2
43468.9 0
0
8 Battery~
219 362 109 0 2 5
0 4 6
0
0 0 880 90
3 0.7
-11 -21 10 -13
2 V3
-8 -31 6 -23
0
0
14 %D %1 %2 DC %V
0
0
0
5

0 1 2 1 2 0
86 0 0 0 0 0 0 0
1 V
8157 0 0
2
43468.9 0
0
8 Battery~
219 298 222 0 2 5
0 5 2
0
0 0 880 0
3 12V
12 -2 33 6
2 V1
16 -12 30 -4
0
0
14 %D %1 %2 DC %V
0
0
0
5

0 1 2 1 2 0
86 0 0 0 0 0 0 0
1 V
5572 0 0
2
43468.9 0
0
9 Resistor~
219 561 169 0 2 5
0 2 3
0
0 0 880 90
8 5.6k Ohm
-13 0 43 8
2 R1
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 0 0 0 0
1 R
8901 0 0
2
43468.9 0
0
8
1 0 0 0 0 0 0 3 0 0 8 2
373 275
373 242
4 0 2 0 0 4096 0 1 0 0 8 2
655 195
561 195
1 0 3 0 0 4096 0 1 0 0 7 2
655 145
561 145
4 1 4 0 0 4224 0 2 5 0 0 4
299 126
336 126
336 106
352 106
1 1 5 0 0 4240 0 6 2 0 0 3
298 209
298 176
299 176
2 1 6 0 0 4224 0 5 4 0 0 2
376 106
431 106
2 2 3 0 0 4224 0 4 7 0 0 3
455 106
561 106
561 151
2 1 2 0 0 8320 0 6 7 0 0 4
298 233
298 242
561 242
561 187
0
0
2049 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
